package cpu_constants is
  constant word_width : integer := 7;
end package;
