library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;

entity control_unit is
  port (Clock       : in std_logic;
        reset       : in std_logic;
        w         : out std_logic);
end entity;

architecture control_unit_arch of control_unit is

begin

end architecture;
